PSpice application example using MC33363 and TL431
.TRAN 50n 10.05m 10m 100n UIC
.OPTIONS abstol=1U itl5=0
.OPTIONS gmin=10n reltol=0.01 vntol=1M
.LIB MC33363.LIB
.PROBE
.PARAM RDSON=15 	; change this parameter if you use 363A or 363B
R4 22 23 2.8k
R1 0 1 15k
C1 0 2 820p
Vin VHT 0 DC=320
X2 8 Prim 14 26 XFMR PARAMS: RATIO={-0.065}
L1 8 3 1M
R2 3 Prim 1.2
D1 14 24 DN5818
C2 21 26 220U
R3 22 26 3
X1 16 Aux 0 0 1 2 REF CMP REF 13 0 0 5 MC33363 PARAMS: RDSON={RDSON}
X4 8 Prim 11 0 XFMR PARAMS: RATIO={-0.169}
R5 23 26 2.74k
Lleak Prim 5 10uH
D2 11 18 MUR120
R6 18 Aux 39
V2 VHT 8
V3 VHT 16
X5 7 26 23 TL431
R9 21 22 100m
C4 Aux 0 10U IC=15
R10 4 8 100k
C5 8 4 1nF
X6 19 7 CMP 0 MOC8101
C6 8 15 47P
R11 15 5 2.2K
R12 24 19 220
R15 24 6 20m
C3 6 26 1000U IC=0
R14 CMP REF 2.7k
L2 24 28 5U
C8 7 23 100N IC=4.5
R16 28 22 10m
R17 Aux 13 5.1k
R18 13 0 1k
D4 5 4 MUR160
Rconv 26 0 10Meg
.END
