* PSpice application file for revised CS5323
.TRAN 0.05u 1.10m 1.05m 0.05u UIC
.LIB D:CS5323.LIB
.OPTIONS abstol=1u itl4=500
.OPTIONS gmin=10n reltol=0.01 vntol=1m
.PROBE
Rdummy 131 0 1Meg
D3 14 28 DKEH 
R14 11 10 2.7K
C23 8 32 0.01U
C12 4 3 1N IC=-10
C13 13 34 540U IC=12
R1 14 15 10
C24 9 32 0.01U
R15 7 25 30.1K
D5 14 112 DKEH 
C4 33 25 1.0U
C25 11 0 0.1U IC=3.3
R16 8 16 30.1K
C14 3 0 0.1U IC=2.2
Resr0 34 0 0.04
C26 112 27 1.0U
RLOAD 32 0 41m
C5 14 0 1.0U
R17 9 27 30.1K
R_L2 32 17 0.01M
C27 14 0 1.0U
C16 32 22 4480U IC=1.7
R18 10 0 1.0K
R_L3 32 20 0.01M
R19 14 131 10K
X_U1 25 44 33 1 131 14 23 0 SC1205
C17 15 0 0.01U IC=5
C28 5 32 1.0N
R_L4 32 21 0.01M
C18 28 16 1.0U
V5IN 14 0 DC=5
R6 5 12 7.5K
X_U2 74 4 5 12 7 8 9 6 10 11 0 11 11 0 0 0 18 2 1 15 CS5323
L1 19 13 300N IC=5
C19 14 0 1.0U
X_U3 16 38 28 2 131 14 43 0 SC1205
V12IN 19 0 DC=12
X_U4 27 46 112 18 131 14 51 0 SC1205
L2 25 17 850N
X_Q1 13 44 25 MTD3302
L3 16 20 850N
R9 5 32 1K
X_Q2 25 23 0 MTD3302
L4 27 21 850N
X_Q3 13 38 16 MTD3302
Resr1 22 0 1.5M
X_Q4 16 43 0 MTD3302
RCORE 19 13 1K
X_Q5 13 46 27 MTD3302
R10 4 3 8K
X_Q6 27 51 0 MTD3302
D1 14 33 DKEH 
C10 32 24 30U IC=1.7
R12 74 0 75K
C21 32 0 0.01U
R13 32 6 10K
C22 7 32 0.01U
C11 4 5 2N
Resr2 0 24 0.15
.MODEL DKEH D
.END
