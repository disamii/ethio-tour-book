* PSpice CS5307 application example
.LIB G:CS5307.LIB
.TRAN 100N 450U 400U 50N UIC
.OPTIONS itl1=1000 itl4=100
.OPTIONS gmin=10n reltol=0.01
.OPTIONS ABSTOL=10u VNTOL=10m
.PROBE
C1 5 0 0.01N
V1 18 0 DC=5
R8 0 17 2m
R1 0 1 32.4k
C5 21 23 1.0U
X1 0 1 1 8 9 10 13 7 42 38 6 5 20 0 0 2 0 0 2 400 300 200 100 24 CS5307
V2 24 0 DC=12
RLOAD 0 7 18.75m
D1 18 21 _D4_mod 
D2 18 16 _D4_mod 
D7 18 22 _D4_mod 
C11 7 17 4480U
R7 13 12 24.9K
C8 13 7 0.01U
X_U1 23 25 21 100 18 18 19 0 SC1205
R9 8 23 24.9K
C9 8 7 0.01U
R10 9 27 24.9K
C10 10 7 0.01U
R11 10 15 24.9K
L1 23 32 820N
X_Q1 4 25 23 mtd3302
C14 9 7 0.01U
X_Q2 23 19 0 mtd3302
V3 2 0 DC=3.3
R12 24 20 5k
C15 6 0 1N
R13 7 38 1.94K
R14 42 38 38.5K
L5 24 4 300N
C17 4 43 540U
C16 7 3 30U
Resr2 3 0 0.15
R_L1 32 7 3.3m
C2 14 27 1.0U
X11 27 31 14 200 18 18 29 0 SC1205
X12 4 31 27 mtd3302
X13 27 29 0 mtd3302
D4 18 14 _D4_mod 
C3 15 16 1.0U
X14 15 41 16 300 18 18 36 0 SC1205
X15 4 41 15 mtd3302
X16 15 36 0 mtd3302
R15 43 0 0.14
C4 22 12 1.0U
X17 12 33 22 400 18 18 40 0 SC1205
X18 4 33 12 mtd3302
X19 12 40 0 mtd3302
Rcore 24 4 1k
C6 18 0 1.0U
C7 18 0 1.0U
C12 18 0 1.0U
C13 18 0 1.0U
L2 27 26 820N
R_L2 26 7 3.3m
L3 15 28 820N
R_L3 28 7 3.3m
L4 12 39 820N
R_L4 39 7 3.3m
.MODEL _D4_mod D (RS=0.78 N=1.95 IS=7.075E-9 
+ CJO=4P TT=7.2N M=.4 VJ=.657 BV=100 IBV=100U)
.END
