MC44608 PSpice demo circuit in a three output 100W SMPS
.LIB MC44608.LIB
.TRAN 1U 100U
.AC DEC 100 1 100k
.PROBE
.PARAM FSW=75k			; switching frequency
.PARAM LP=180u			; primary inductance
.PARAM RATIO8V=0.071	; XFMR ratio for 8V output
.PARAM RATIO18V=0.2		; XFMR ratio for 18V output
.PARAM RATIO112V=1		; XFMR ratio for 112V output
X1 9 9 2 0 6 20 MC44608 PARAMS: Lp={LP} Fs={FSW}
C1 Vout 4 47uF
R1 4 0 400m
V2 Vout 12
R7 2 0 10k
V1 20 0 DC=370	; DC Input voltage, AC statement sweeps audio
R3 8 2 100
Vdc 8 0 DC=5.26 AC=1 ; Duty-cycle set point and AC stimulus
R2 12 0 180	; 112V output
X6 6 0 19 0 XFMR1 PARAMS: RATIO={RATIO112V}
C4 7 0 1mF
R9 V8 7 500m
V5 V8 1
R10 1 0 8	; 8V output
X4 6 0 16 0 XFMR1 PARAMS: RATIO={RATIO8V}
D4 19 Vout MR854
C5 V18 21 1mF
R11 21 0 500m
V6 V18 22	; 18V output
R12 22 0 18
X7 6 0 23 0 XFMR1 PARAMS: RATIO={RATIO18V}
D6 23 V18 MR852
D7 16 V8 MR852
.MODEL MR854 D BV=400 CJO=124P IBV=100N IS=3.91N M=.333
+ N=1.67 RS=14.6M TT=520N VJ=.75
.MODEL MR852 D BV=200 CJO=124P IBV=100N IS=3.91N M=.333
+ N=1.67 RS=14.6M TT=520N VJ=.75
.END
