* CS5322 Application example
.TRAN 100n 1020u 1000u 50N UIC
.OPTIONS itl4=1000
.PROBE
.LIB D:CS5322.LIB
Rdummy 21 0 10Meg
R14 27 25 4.32K
RESR_C3 9 0 4.3M
C2 8 11 6560U
R15 27 0 1K
C3 3 9 2040U IC=5
R16 6 1 2K
C5 12 0 0.01U
R3 8 0 45.7M
R_L1 4 8 1.25M
C6 19 0 1N
R_L2 5 8 1.25M
C7 19 22 1N
R5 0 11 1.5M
C8 8 23 0.01U
C9 8 24 0.01U
L1 10 4 470N
R8 0 17 61.9K
L2 2 5 470N
R9 22 18 25.5K
L3 6 3 300N
X1 19 22 18 24 23 21 1 0 25 0 25 0 27 25 15 13 0 14 6 12 0
+ 15 20 0 16 6 6 17 CS5322
R10 22 8 7.5K
RCORE 6 3 1K
X2 3 20 10 MTD3302
R11 8 21 12.7K
V1 6 0 DC=5V
X3 10 16 0 MTD3302
C10 25 0 0.1U
R12 23 2 25.5K
V2 15 0 DC=12
RESR_C1 7 0 37.5M
X4 3 13 2 MTD3302
R13 24 10 25.5K
C1 8 7 120U
X5 2 14 0 MTD3302
.END
